library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity Ascen is

    
end Ascen;

architecture Behavioral of Ascen is

begin


end Behavioral;
